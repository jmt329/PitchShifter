module delta_rom (clock, address, delta_out);
   input clock;
   input [9:0] address;
   output [31:0] delta_out;
   reg [31:0]    delta_out;
   always@(posedge clock)
     begin
        case(address)
          10'd0: delta_out   = 32'b00010000000000000000000000000000;
          10'd1: delta_out   = 32'b00010000001000000000000000000000;
          10'd2: delta_out   = 32'b00010000010000000000000000000000;
          10'd3: delta_out   = 32'b00010000011000000000000000000000;
          10'd4: delta_out   = 32'b00010000100000000000000000000000;
          10'd5: delta_out   = 32'b00010000101000000000000000000000;
          10'd6: delta_out   = 32'b00010000110000000000000000000000;
          10'd7: delta_out   = 32'b00010000111000000000000000000000;
          10'd8: delta_out   = 32'b00010001000000000000000000000000;
          10'd9: delta_out   = 32'b00010001001000000000000000000000;
          10'd10: delta_out  = 32'b00010001010000000000000000000000;
          10'd11: delta_out  = 32'b00010001011000000000000000000000;
          10'd12: delta_out  = 32'b00010001100000000000000000000000;
          10'd13: delta_out  = 32'b00010001101000000000000000000000;
          10'd14: delta_out  = 32'b00010001110000000000000000000000;
          10'd15: delta_out  = 32'b00010001111000000000000000000000;
          10'd16: delta_out  = 32'b00010010000000000000000000000000;
          10'd17: delta_out  = 32'b00010010001000000000000000000000;
          10'd18: delta_out  = 32'b00010010010000000000000000000000;
          10'd19: delta_out  = 32'b00010010011000000000000000000000;
          10'd20: delta_out  = 32'b00010010100000000000000000000000;
          10'd21: delta_out  = 32'b00010010101000000000000000000000;
          10'd22: delta_out  = 32'b00010010110000000000000000000000;
          10'd23: delta_out  = 32'b00010010111000000000000000000000;
          10'd24: delta_out  = 32'b00010011000000000000000000000000;
          10'd25: delta_out  = 32'b00010011001000000000000000000000;
          10'd26: delta_out  = 32'b00010011010000000000000000000000;
          10'd27: delta_out  = 32'b00010011011000000000000000000000;
          10'd28: delta_out  = 32'b00010011100000000000000000000000;
          10'd29: delta_out  = 32'b00010011101000000000000000000000;
          10'd30: delta_out  = 32'b00010011110000000000000000000000;
          10'd31: delta_out  = 32'b00010011111000000000000000000000;
          10'd32: delta_out  = 32'b00010100000000000000000000000000;
          10'd33: delta_out  = 32'b00010100001000000000000000000000;
          10'd34: delta_out  = 32'b00010100010000000000000000000000;
          10'd35: delta_out  = 32'b00010100011000000000000000000000;
          10'd36: delta_out  = 32'b00010100100000000000000000000000;
          10'd37: delta_out  = 32'b00010100101000000000000000000000;
          10'd38: delta_out  = 32'b00010100110000000000000000000000;
          10'd39: delta_out  = 32'b00010100111000000000000000000000;
          10'd40: delta_out  = 32'b00010101000000000000000000000000;
          10'd41: delta_out  = 32'b00010101001000000000000000000000;
          10'd42: delta_out  = 32'b00010101010000000000000000000000;
          10'd43: delta_out  = 32'b00010101011000000000000000000000;
          10'd44: delta_out  = 32'b00010101100000000000000000000000;
          10'd45: delta_out  = 32'b00010101101000000000000000000000;
          10'd46: delta_out  = 32'b00010101110000000000000000000000;
          10'd47: delta_out  = 32'b00010101111000000000000000000000;
          10'd48: delta_out  = 32'b00010110000000000000000000000000;
          10'd49: delta_out  = 32'b00010110001000000000000000000000;
          10'd50: delta_out  = 32'b00010110010000000000000000000000;
          10'd51: delta_out  = 32'b00010110011000000000000000000000;
          10'd52: delta_out  = 32'b00010110100000000000000000000000;
          10'd53: delta_out  = 32'b00010110101000000000000000000000;
          10'd54: delta_out  = 32'b00010110110000000000000000000000;
          10'd55: delta_out  = 32'b00010110111000000000000000000000;
          10'd56: delta_out  = 32'b00010111000000000000000000000000;
          10'd57: delta_out  = 32'b00010111001000000000000000000000;
          10'd58: delta_out  = 32'b00010111010000000000000000000000;
          10'd59: delta_out  = 32'b00010111011000000000000000000000;
          10'd60: delta_out  = 32'b00010111100000000000000000000000;
          10'd61: delta_out  = 32'b00010111101000000000000000000000;
          10'd62: delta_out  = 32'b00010111110000000000000000000000;
          10'd63: delta_out  = 32'b00010111111000000000000000000000;
          10'd64: delta_out  = 32'b00011000000000000000000000000000;
          10'd65: delta_out  = 32'b00011000001000000000000000000000;
          10'd66: delta_out  = 32'b00011000010000000000000000000000;
          10'd67: delta_out  = 32'b00011000011000000000000000000000;
          10'd68: delta_out  = 32'b00011000100000000000000000000000;
          10'd69: delta_out  = 32'b00011000101000000000000000000000;
          10'd70: delta_out  = 32'b00011000110000000000000000000000;
          10'd71: delta_out  = 32'b00011000111000000000000000000000;
          10'd72: delta_out  = 32'b00011001000000000000000000000000;
          10'd73: delta_out  = 32'b00011001001000000000000000000000;
          10'd74: delta_out  = 32'b00011001010000000000000000000000;
          10'd75: delta_out  = 32'b00011001011000000000000000000000;
          10'd76: delta_out  = 32'b00011001100000000000000000000000;
          10'd77: delta_out  = 32'b00011001101000000000000000000000;
          10'd78: delta_out  = 32'b00011001110000000000000000000000;
          10'd79: delta_out  = 32'b00011001111000000000000000000000;
          10'd80: delta_out  = 32'b00011010000000000000000000000000;
          10'd81: delta_out  = 32'b00011010001000000000000000000000;
          10'd82: delta_out  = 32'b00011010010000000000000000000000;
          10'd83: delta_out  = 32'b00011010011000000000000000000000;
          10'd84: delta_out  = 32'b00011010100000000000000000000000;
          10'd85: delta_out  = 32'b00011010101000000000000000000000;
          10'd86: delta_out  = 32'b00011010110000000000000000000000;
          10'd87: delta_out  = 32'b00011010111000000000000000000000;
          10'd88: delta_out  = 32'b00011011000000000000000000000000;
          10'd89: delta_out  = 32'b00011011001000000000000000000000;
          10'd90: delta_out  = 32'b00011011010000000000000000000000;
          10'd91: delta_out  = 32'b00011011011000000000000000000000;
          10'd92: delta_out  = 32'b00011011100000000000000000000000;
          10'd93: delta_out  = 32'b00011011101000000000000000000000;
          10'd94: delta_out  = 32'b00011011110000000000000000000000;
          10'd95: delta_out  = 32'b00011011111000000000000000000000;
          10'd96: delta_out  = 32'b00011100000000000000000000000000;
          10'd97: delta_out  = 32'b00011100001000000000000000000000;
          10'd98: delta_out  = 32'b00011100010000000000000000000000;
          10'd99: delta_out  = 32'b00011100011000000000000000000000;
          10'd100: delta_out = 32'b00011100100000000000000000000000;
          10'd101: delta_out = 32'b00011100101000000000000000000000;
          10'd102: delta_out = 32'b00011100110000000000000000000000;
          10'd103: delta_out = 32'b00011100111000000000000000000000;
          10'd104: delta_out = 32'b00011101000000000000000000000000;
          10'd105: delta_out = 32'b00011101001000000000000000000000;
          10'd106: delta_out = 32'b00011101010000000000000000000000;
          10'd107: delta_out = 32'b00011101011000000000000000000000;
          10'd108: delta_out = 32'b00011101100000000000000000000000;
          10'd109: delta_out = 32'b00011101101000000000000000000000;
          10'd110: delta_out = 32'b00011101110000000000000000000000;
          10'd111: delta_out = 32'b00011101111000000000000000000000;
          10'd112: delta_out = 32'b00011110000000000000000000000000;
          10'd113: delta_out = 32'b00011110001000000000000000000000;
          10'd114: delta_out = 32'b00011110010000000000000000000000;
          10'd115: delta_out = 32'b00011110011000000000000000000000;
          10'd116: delta_out = 32'b00011110100000000000000000000000;
          10'd117: delta_out = 32'b00011110101000000000000000000000;
          10'd118: delta_out = 32'b00011110110000000000000000000000;
          10'd119: delta_out = 32'b00011110111000000000000000000000;
          10'd120: delta_out = 32'b00011111000000000000000000000000;
          10'd121: delta_out = 32'b00011111001000000000000000000000;
          10'd122: delta_out = 32'b00011111010000000000000000000000;
          10'd123: delta_out = 32'b00011111011000000000000000000000;
          10'd124: delta_out = 32'b00011111100000000000000000000000;
          10'd125: delta_out = 32'b00011111101000000000000000000000;
          10'd126: delta_out = 32'b00011111110000000000000000000000;
          10'd127: delta_out = 32'b00011111111000000000000000000000;
          10'd128: delta_out = 32'b00100000000000000000000000000000;
          10'd129: delta_out = 32'b00100000001000000000000000000000;
          10'd130: delta_out = 32'b00100000010000000000000000000000;
          10'd131: delta_out = 32'b00100000011000000000000000000000;
          10'd132: delta_out = 32'b00100000100000000000000000000000;
          10'd133: delta_out = 32'b00100000101000000000000000000000;
          10'd134: delta_out = 32'b00100000110000000000000000000000;
          10'd135: delta_out = 32'b00100000111000000000000000000000;
          10'd136: delta_out = 32'b00100001000000000000000000000000;
          10'd137: delta_out = 32'b00100001001000000000000000000000;
          10'd138: delta_out = 32'b00100001010000000000000000000000;
          10'd139: delta_out = 32'b00100001011000000000000000000000;
          10'd140: delta_out = 32'b00100001100000000000000000000000;
          10'd141: delta_out = 32'b00100001101000000000000000000000;
          10'd142: delta_out = 32'b00100001110000000000000000000000;
          10'd143: delta_out = 32'b00100001111000000000000000000000;
          10'd144: delta_out = 32'b00100010000000000000000000000000;
          10'd145: delta_out = 32'b00100010001000000000000000000000;
          10'd146: delta_out = 32'b00100010010000000000000000000000;
          10'd147: delta_out = 32'b00100010011000000000000000000000;
          10'd148: delta_out = 32'b00100010100000000000000000000000;
          10'd149: delta_out = 32'b00100010101000000000000000000000;
          10'd150: delta_out = 32'b00100010110000000000000000000000;
          10'd151: delta_out = 32'b00100010111000000000000000000000;
          10'd152: delta_out = 32'b00100011000000000000000000000000;
          10'd153: delta_out = 32'b00100011001000000000000000000000;
          10'd154: delta_out = 32'b00100011010000000000000000000000;
          10'd155: delta_out = 32'b00100011011000000000000000000000;
          10'd156: delta_out = 32'b00100011100000000000000000000000;
          10'd157: delta_out = 32'b00100011101000000000000000000000;
          10'd158: delta_out = 32'b00100011110000000000000000000000;
          10'd159: delta_out = 32'b00100011111000000000000000000000;
          10'd160: delta_out = 32'b00100100000000000000000000000000;
          10'd161: delta_out = 32'b00100100001000000000000000000000;
          10'd162: delta_out = 32'b00100100010000000000000000000000;
          10'd163: delta_out = 32'b00100100011000000000000000000000;
          10'd164: delta_out = 32'b00100100100000000000000000000000;
          10'd165: delta_out = 32'b00100100101000000000000000000000;
          10'd166: delta_out = 32'b00100100110000000000000000000000;
          10'd167: delta_out = 32'b00100100111000000000000000000000;
          10'd168: delta_out = 32'b00100101000000000000000000000000;
          10'd169: delta_out = 32'b00100101001000000000000000000000;
          10'd170: delta_out = 32'b00100101010000000000000000000000;
          10'd171: delta_out = 32'b00100101011000000000000000000000;
          10'd172: delta_out = 32'b00100101100000000000000000000000;
          10'd173: delta_out = 32'b00100101101000000000000000000000;
          10'd174: delta_out = 32'b00100101110000000000000000000000;
          10'd175: delta_out = 32'b00100101111000000000000000000000;
          10'd176: delta_out = 32'b00100110000000000000000000000000;
          10'd177: delta_out = 32'b00100110001000000000000000000000;
          10'd178: delta_out = 32'b00100110010000000000000000000000;
          10'd179: delta_out = 32'b00100110011000000000000000000000;
          10'd180: delta_out = 32'b00100110100000000000000000000000;
          10'd181: delta_out = 32'b00100110101000000000000000000000;
          10'd182: delta_out = 32'b00100110110000000000000000000000;
          10'd183: delta_out = 32'b00100110111000000000000000000000;
          10'd184: delta_out = 32'b00100111000000000000000000000000;
          10'd185: delta_out = 32'b00100111001000000000000000000000;
          10'd186: delta_out = 32'b00100111010000000000000000000000;
          10'd187: delta_out = 32'b00100111011000000000000000000000;
          10'd188: delta_out = 32'b00100111100000000000000000000000;
          10'd189: delta_out = 32'b00100111101000000000000000000000;
          10'd190: delta_out = 32'b00100111110000000000000000000000;
          10'd191: delta_out = 32'b00100111111000000000000000000000;
          10'd192: delta_out = 32'b00101000000000000000000000000000;
          10'd193: delta_out = 32'b00101000001000000000000000000000;
          10'd194: delta_out = 32'b00101000010000000000000000000000;
          10'd195: delta_out = 32'b00101000011000000000000000000000;
          10'd196: delta_out = 32'b00101000100000000000000000000000;
          10'd197: delta_out = 32'b00101000101000000000000000000000;
          10'd198: delta_out = 32'b00101000110000000000000000000000;
          10'd199: delta_out = 32'b00101000111000000000000000000000;
          10'd200: delta_out = 32'b00101001000000000000000000000000;
          10'd201: delta_out = 32'b00101001001000000000000000000000;
          10'd202: delta_out = 32'b00101001010000000000000000000000;
          10'd203: delta_out = 32'b00101001011000000000000000000000;
          10'd204: delta_out = 32'b00101001100000000000000000000000;
          10'd205: delta_out = 32'b00101001101000000000000000000000;
          10'd206: delta_out = 32'b00101001110000000000000000000000;
          10'd207: delta_out = 32'b00101001111000000000000000000000;
          10'd208: delta_out = 32'b00101010000000000000000000000000;
          10'd209: delta_out = 32'b00101010001000000000000000000000;
          10'd210: delta_out = 32'b00101010010000000000000000000000;
          10'd211: delta_out = 32'b00101010011000000000000000000000;
          10'd212: delta_out = 32'b00101010100000000000000000000000;
          10'd213: delta_out = 32'b00101010101000000000000000000000;
          10'd214: delta_out = 32'b00101010110000000000000000000000;
          10'd215: delta_out = 32'b00101010111000000000000000000000;
          10'd216: delta_out = 32'b00101011000000000000000000000000;
          10'd217: delta_out = 32'b00101011001000000000000000000000;
          10'd218: delta_out = 32'b00101011010000000000000000000000;
          10'd219: delta_out = 32'b00101011011000000000000000000000;
          10'd220: delta_out = 32'b00101011100000000000000000000000;
          10'd221: delta_out = 32'b00101011101000000000000000000000;
          10'd222: delta_out = 32'b00101011110000000000000000000000;
          10'd223: delta_out = 32'b00101011111000000000000000000000;
          10'd224: delta_out = 32'b00101100000000000000000000000000;
          10'd225: delta_out = 32'b00101100001000000000000000000000;
          10'd226: delta_out = 32'b00101100010000000000000000000000;
          10'd227: delta_out = 32'b00101100011000000000000000000000;
          10'd228: delta_out = 32'b00101100100000000000000000000000;
          10'd229: delta_out = 32'b00101100101000000000000000000000;
          10'd230: delta_out = 32'b00101100110000000000000000000000;
          10'd231: delta_out = 32'b00101100111000000000000000000000;
          10'd232: delta_out = 32'b00101101000000000000000000000000;
          10'd233: delta_out = 32'b00101101001000000000000000000000;
          10'd234: delta_out = 32'b00101101010000000000000000000000;
          10'd235: delta_out = 32'b00101101011000000000000000000000;
          10'd236: delta_out = 32'b00101101100000000000000000000000;
          10'd237: delta_out = 32'b00101101101000000000000000000000;
          10'd238: delta_out = 32'b00101101110000000000000000000000;
          10'd239: delta_out = 32'b00101101111000000000000000000000;
          10'd240: delta_out = 32'b00101110000000000000000000000000;
          10'd241: delta_out = 32'b00101110001000000000000000000000;
          10'd242: delta_out = 32'b00101110010000000000000000000000;
          10'd243: delta_out = 32'b00101110011000000000000000000000;
          10'd244: delta_out = 32'b00101110100000000000000000000000;
          10'd245: delta_out = 32'b00101110101000000000000000000000;
          10'd246: delta_out = 32'b00101110110000000000000000000000;
          10'd247: delta_out = 32'b00101110111000000000000000000000;
          10'd248: delta_out = 32'b00101111000000000000000000000000;
          10'd249: delta_out = 32'b00101111001000000000000000000000;
          10'd250: delta_out = 32'b00101111010000000000000000000000;
          10'd251: delta_out = 32'b00101111011000000000000000000000;
          10'd252: delta_out = 32'b00101111100000000000000000000000;
          10'd253: delta_out = 32'b00101111101000000000000000000000;
          10'd254: delta_out = 32'b00101111110000000000000000000000;
          10'd255: delta_out = 32'b00101111111000000000000000000000;
          10'd256: delta_out = 32'b00110000000000000000000000000000;
          10'd257: delta_out = 32'b00101111111000000000000000000000;
          10'd258: delta_out = 32'b00101111110000000000000000000000;
          10'd259: delta_out = 32'b00101111101000000000000000000000;
          10'd260: delta_out = 32'b00101111100000000000000000000000;
          10'd261: delta_out = 32'b00101111011000000000000000000000;
          10'd262: delta_out = 32'b00101111010000000000000000000000;
          10'd263: delta_out = 32'b00101111001000000000000000000000;
          10'd264: delta_out = 32'b00101111000000000000000000000000;
          10'd265: delta_out = 32'b00101110111000000000000000000000;
          10'd266: delta_out = 32'b00101110110000000000000000000000;
          10'd267: delta_out = 32'b00101110101000000000000000000000;
          10'd268: delta_out = 32'b00101110100000000000000000000000;
          10'd269: delta_out = 32'b00101110011000000000000000000000;
          10'd270: delta_out = 32'b00101110010000000000000000000000;
          10'd271: delta_out = 32'b00101110001000000000000000000000;
          10'd272: delta_out = 32'b00101110000000000000000000000000;
          10'd273: delta_out = 32'b00101101111000000000000000000000;
          10'd274: delta_out = 32'b00101101110000000000000000000000;
          10'd275: delta_out = 32'b00101101101000000000000000000000;
          10'd276: delta_out = 32'b00101101100000000000000000000000;
          10'd277: delta_out = 32'b00101101011000000000000000000000;
          10'd278: delta_out = 32'b00101101010000000000000000000000;
          10'd279: delta_out = 32'b00101101001000000000000000000000;
          10'd280: delta_out = 32'b00101101000000000000000000000000;
          10'd281: delta_out = 32'b00101100111000000000000000000000;
          10'd282: delta_out = 32'b00101100110000000000000000000000;
          10'd283: delta_out = 32'b00101100101000000000000000000000;
          10'd284: delta_out = 32'b00101100100000000000000000000000;
          10'd285: delta_out = 32'b00101100011000000000000000000000;
          10'd286: delta_out = 32'b00101100010000000000000000000000;
          10'd287: delta_out = 32'b00101100001000000000000000000000;
          10'd288: delta_out = 32'b00101100000000000000000000000000;
          10'd289: delta_out = 32'b00101011111000000000000000000000;
          10'd290: delta_out = 32'b00101011110000000000000000000000;
          10'd291: delta_out = 32'b00101011101000000000000000000000;
          10'd292: delta_out = 32'b00101011100000000000000000000000;
          10'd293: delta_out = 32'b00101011011000000000000000000000;
          10'd294: delta_out = 32'b00101011010000000000000000000000;
          10'd295: delta_out = 32'b00101011001000000000000000000000;
          10'd296: delta_out = 32'b00101011000000000000000000000000;
          10'd297: delta_out = 32'b00101010111000000000000000000000;
          10'd298: delta_out = 32'b00101010110000000000000000000000;
          10'd299: delta_out = 32'b00101010101000000000000000000000;
          10'd300: delta_out = 32'b00101010100000000000000000000000;
          10'd301: delta_out = 32'b00101010011000000000000000000000;
          10'd302: delta_out = 32'b00101010010000000000000000000000;
          10'd303: delta_out = 32'b00101010001000000000000000000000;
          10'd304: delta_out = 32'b00101010000000000000000000000000;
          10'd305: delta_out = 32'b00101001111000000000000000000000;
          10'd306: delta_out = 32'b00101001110000000000000000000000;
          10'd307: delta_out = 32'b00101001101000000000000000000000;
          10'd308: delta_out = 32'b00101001100000000000000000000000;
          10'd309: delta_out = 32'b00101001011000000000000000000000;
          10'd310: delta_out = 32'b00101001010000000000000000000000;
          10'd311: delta_out = 32'b00101001001000000000000000000000;
          10'd312: delta_out = 32'b00101001000000000000000000000000;
          10'd313: delta_out = 32'b00101000111000000000000000000000;
          10'd314: delta_out = 32'b00101000110000000000000000000000;
          10'd315: delta_out = 32'b00101000101000000000000000000000;
          10'd316: delta_out = 32'b00101000100000000000000000000000;
          10'd317: delta_out = 32'b00101000011000000000000000000000;
          10'd318: delta_out = 32'b00101000010000000000000000000000;
          10'd319: delta_out = 32'b00101000001000000000000000000000;
          10'd320: delta_out = 32'b00101000000000000000000000000000;
          10'd321: delta_out = 32'b00100111111000000000000000000000;
          10'd322: delta_out = 32'b00100111110000000000000000000000;
          10'd323: delta_out = 32'b00100111101000000000000000000000;
          10'd324: delta_out = 32'b00100111100000000000000000000000;
          10'd325: delta_out = 32'b00100111011000000000000000000000;
          10'd326: delta_out = 32'b00100111010000000000000000000000;
          10'd327: delta_out = 32'b00100111001000000000000000000000;
          10'd328: delta_out = 32'b00100111000000000000000000000000;
          10'd329: delta_out = 32'b00100110111000000000000000000000;
          10'd330: delta_out = 32'b00100110110000000000000000000000;
          10'd331: delta_out = 32'b00100110101000000000000000000000;
          10'd332: delta_out = 32'b00100110100000000000000000000000;
          10'd333: delta_out = 32'b00100110011000000000000000000000;
          10'd334: delta_out = 32'b00100110010000000000000000000000;
          10'd335: delta_out = 32'b00100110001000000000000000000000;
          10'd336: delta_out = 32'b00100110000000000000000000000000;
          10'd337: delta_out = 32'b00100101111000000000000000000000;
          10'd338: delta_out = 32'b00100101110000000000000000000000;
          10'd339: delta_out = 32'b00100101101000000000000000000000;
          10'd340: delta_out = 32'b00100101100000000000000000000000;
          10'd341: delta_out = 32'b00100101011000000000000000000000;
          10'd342: delta_out = 32'b00100101010000000000000000000000;
          10'd343: delta_out = 32'b00100101001000000000000000000000;
          10'd344: delta_out = 32'b00100101000000000000000000000000;
          10'd345: delta_out = 32'b00100100111000000000000000000000;
          10'd346: delta_out = 32'b00100100110000000000000000000000;
          10'd347: delta_out = 32'b00100100101000000000000000000000;
          10'd348: delta_out = 32'b00100100100000000000000000000000;
          10'd349: delta_out = 32'b00100100011000000000000000000000;
          10'd350: delta_out = 32'b00100100010000000000000000000000;
          10'd351: delta_out = 32'b00100100001000000000000000000000;
          10'd352: delta_out = 32'b00100100000000000000000000000000;
          10'd353: delta_out = 32'b00100011111000000000000000000000;
          10'd354: delta_out = 32'b00100011110000000000000000000000;
          10'd355: delta_out = 32'b00100011101000000000000000000000;
          10'd356: delta_out = 32'b00100011100000000000000000000000;
          10'd357: delta_out = 32'b00100011011000000000000000000000;
          10'd358: delta_out = 32'b00100011010000000000000000000000;
          10'd359: delta_out = 32'b00100011001000000000000000000000;
          10'd360: delta_out = 32'b00100011000000000000000000000000;
          10'd361: delta_out = 32'b00100010111000000000000000000000;
          10'd362: delta_out = 32'b00100010110000000000000000000000;
          10'd363: delta_out = 32'b00100010101000000000000000000000;
          10'd364: delta_out = 32'b00100010100000000000000000000000;
          10'd365: delta_out = 32'b00100010011000000000000000000000;
          10'd366: delta_out = 32'b00100010010000000000000000000000;
          10'd367: delta_out = 32'b00100010001000000000000000000000;
          10'd368: delta_out = 32'b00100010000000000000000000000000;
          10'd369: delta_out = 32'b00100001111000000000000000000000;
          10'd370: delta_out = 32'b00100001110000000000000000000000;
          10'd371: delta_out = 32'b00100001101000000000000000000000;
          10'd372: delta_out = 32'b00100001100000000000000000000000;
          10'd373: delta_out = 32'b00100001011000000000000000000000;
          10'd374: delta_out = 32'b00100001010000000000000000000000;
          10'd375: delta_out = 32'b00100001001000000000000000000000;
          10'd376: delta_out = 32'b00100001000000000000000000000000;
          10'd377: delta_out = 32'b00100000111000000000000000000000;
          10'd378: delta_out = 32'b00100000110000000000000000000000;
          10'd379: delta_out = 32'b00100000101000000000000000000000;
          10'd380: delta_out = 32'b00100000100000000000000000000000;
          10'd381: delta_out = 32'b00100000011000000000000000000000;
          10'd382: delta_out = 32'b00100000010000000000000000000000;
          10'd383: delta_out = 32'b00100000001000000000000000000000;
          10'd384: delta_out = 32'b00100000000000000000000000000000;
          10'd385: delta_out = 32'b00011111111000000000000000000000;
          10'd386: delta_out = 32'b00011111110000000000000000000000;
          10'd387: delta_out = 32'b00011111101000000000000000000000;
          10'd388: delta_out = 32'b00011111100000000000000000000000;
          10'd389: delta_out = 32'b00011111011000000000000000000000;
          10'd390: delta_out = 32'b00011111010000000000000000000000;
          10'd391: delta_out = 32'b00011111001000000000000000000000;
          10'd392: delta_out = 32'b00011111000000000000000000000000;
          10'd393: delta_out = 32'b00011110111000000000000000000000;
          10'd394: delta_out = 32'b00011110110000000000000000000000;
          10'd395: delta_out = 32'b00011110101000000000000000000000;
          10'd396: delta_out = 32'b00011110100000000000000000000000;
          10'd397: delta_out = 32'b00011110011000000000000000000000;
          10'd398: delta_out = 32'b00011110010000000000000000000000;
          10'd399: delta_out = 32'b00011110001000000000000000000000;
          10'd400: delta_out = 32'b00011110000000000000000000000000;
          10'd401: delta_out = 32'b00011101111000000000000000000000;
          10'd402: delta_out = 32'b00011101110000000000000000000000;
          10'd403: delta_out = 32'b00011101101000000000000000000000;
          10'd404: delta_out = 32'b00011101100000000000000000000000;
          10'd405: delta_out = 32'b00011101011000000000000000000000;
          10'd406: delta_out = 32'b00011101010000000000000000000000;
          10'd407: delta_out = 32'b00011101001000000000000000000000;
          10'd408: delta_out = 32'b00011101000000000000000000000000;
          10'd409: delta_out = 32'b00011100111000000000000000000000;
          10'd410: delta_out = 32'b00011100110000000000000000000000;
          10'd411: delta_out = 32'b00011100101000000000000000000000;
          10'd412: delta_out = 32'b00011100100000000000000000000000;
          10'd413: delta_out = 32'b00011100011000000000000000000000;
          10'd414: delta_out = 32'b00011100010000000000000000000000;
          10'd415: delta_out = 32'b00011100001000000000000000000000;
          10'd416: delta_out = 32'b00011100000000000000000000000000;
          10'd417: delta_out = 32'b00011011111000000000000000000000;
          10'd418: delta_out = 32'b00011011110000000000000000000000;
          10'd419: delta_out = 32'b00011011101000000000000000000000;
          10'd420: delta_out = 32'b00011011100000000000000000000000;
          10'd421: delta_out = 32'b00011011011000000000000000000000;
          10'd422: delta_out = 32'b00011011010000000000000000000000;
          10'd423: delta_out = 32'b00011011001000000000000000000000;
          10'd424: delta_out = 32'b00011011000000000000000000000000;
          10'd425: delta_out = 32'b00011010111000000000000000000000;
          10'd426: delta_out = 32'b00011010110000000000000000000000;
          10'd427: delta_out = 32'b00011010101000000000000000000000;
          10'd428: delta_out = 32'b00011010100000000000000000000000;
          10'd429: delta_out = 32'b00011010011000000000000000000000;
          10'd430: delta_out = 32'b00011010010000000000000000000000;
          10'd431: delta_out = 32'b00011010001000000000000000000000;
          10'd432: delta_out = 32'b00011010000000000000000000000000;
          10'd433: delta_out = 32'b00011001111000000000000000000000;
          10'd434: delta_out = 32'b00011001110000000000000000000000;
          10'd435: delta_out = 32'b00011001101000000000000000000000;
          10'd436: delta_out = 32'b00011001100000000000000000000000;
          10'd437: delta_out = 32'b00011001011000000000000000000000;
          10'd438: delta_out = 32'b00011001010000000000000000000000;
          10'd439: delta_out = 32'b00011001001000000000000000000000;
          10'd440: delta_out = 32'b00011001000000000000000000000000;
          10'd441: delta_out = 32'b00011000111000000000000000000000;
          10'd442: delta_out = 32'b00011000110000000000000000000000;
          10'd443: delta_out = 32'b00011000101000000000000000000000;
          10'd444: delta_out = 32'b00011000100000000000000000000000;
          10'd445: delta_out = 32'b00011000011000000000000000000000;
          10'd446: delta_out = 32'b00011000010000000000000000000000;
          10'd447: delta_out = 32'b00011000001000000000000000000000;
          10'd448: delta_out = 32'b00011000000000000000000000000000;
          10'd449: delta_out = 32'b00010111111000000000000000000000;
          10'd450: delta_out = 32'b00010111110000000000000000000000;
          10'd451: delta_out = 32'b00010111101000000000000000000000;
          10'd452: delta_out = 32'b00010111100000000000000000000000;
          10'd453: delta_out = 32'b00010111011000000000000000000000;
          10'd454: delta_out = 32'b00010111010000000000000000000000;
          10'd455: delta_out = 32'b00010111001000000000000000000000;
          10'd456: delta_out = 32'b00010111000000000000000000000000;
          10'd457: delta_out = 32'b00010110111000000000000000000000;
          10'd458: delta_out = 32'b00010110110000000000000000000000;
          10'd459: delta_out = 32'b00010110101000000000000000000000;
          10'd460: delta_out = 32'b00010110100000000000000000000000;
          10'd461: delta_out = 32'b00010110011000000000000000000000;
          10'd462: delta_out = 32'b00010110010000000000000000000000;
          10'd463: delta_out = 32'b00010110001000000000000000000000;
          10'd464: delta_out = 32'b00010110000000000000000000000000;
          10'd465: delta_out = 32'b00010101111000000000000000000000;
          10'd466: delta_out = 32'b00010101110000000000000000000000;
          10'd467: delta_out = 32'b00010101101000000000000000000000;
          10'd468: delta_out = 32'b00010101100000000000000000000000;
          10'd469: delta_out = 32'b00010101011000000000000000000000;
          10'd470: delta_out = 32'b00010101010000000000000000000000;
          10'd471: delta_out = 32'b00010101001000000000000000000000;
          10'd472: delta_out = 32'b00010101000000000000000000000000;
          10'd473: delta_out = 32'b00010100111000000000000000000000;
          10'd474: delta_out = 32'b00010100110000000000000000000000;
          10'd475: delta_out = 32'b00010100101000000000000000000000;
          10'd476: delta_out = 32'b00010100100000000000000000000000;
          10'd477: delta_out = 32'b00010100011000000000000000000000;
          10'd478: delta_out = 32'b00010100010000000000000000000000;
          10'd479: delta_out = 32'b00010100001000000000000000000000;
          10'd480: delta_out = 32'b00010100000000000000000000000000;
          10'd481: delta_out = 32'b00010011111000000000000000000000;
          10'd482: delta_out = 32'b00010011110000000000000000000000;
          10'd483: delta_out = 32'b00010011101000000000000000000000;
          10'd484: delta_out = 32'b00010011100000000000000000000000;
          10'd485: delta_out = 32'b00010011011000000000000000000000;
          10'd486: delta_out = 32'b00010011010000000000000000000000;
          10'd487: delta_out = 32'b00010011001000000000000000000000;
          10'd488: delta_out = 32'b00010011000000000000000000000000;
          10'd489: delta_out = 32'b00010010111000000000000000000000;
          10'd490: delta_out = 32'b00010010110000000000000000000000;
          10'd491: delta_out = 32'b00010010101000000000000000000000;
          10'd492: delta_out = 32'b00010010100000000000000000000000;
          10'd493: delta_out = 32'b00010010011000000000000000000000;
          10'd494: delta_out = 32'b00010010010000000000000000000000;
          10'd495: delta_out = 32'b00010010001000000000000000000000;
          10'd496: delta_out = 32'b00010010000000000000000000000000;
          10'd497: delta_out = 32'b00010001111000000000000000000000;
          10'd498: delta_out = 32'b00010001110000000000000000000000;
          10'd499: delta_out = 32'b00010001101000000000000000000000;
          10'd500: delta_out = 32'b00010001100000000000000000000000;
          10'd501: delta_out = 32'b00010001011000000000000000000000;
          10'd502: delta_out = 32'b00010001010000000000000000000000;
          10'd503: delta_out = 32'b00010001001000000000000000000000;
          10'd504: delta_out = 32'b00010001000000000000000000000000;
          10'd505: delta_out = 32'b00010000111000000000000000000000;
          10'd506: delta_out = 32'b00010000110000000000000000000000;
          10'd507: delta_out = 32'b00010000101000000000000000000000;
          10'd508: delta_out = 32'b00010000100000000000000000000000;
          10'd509: delta_out = 32'b00010000011000000000000000000000;
          10'd510: delta_out = 32'b00010000010000000000000000000000;
          10'd511: delta_out = 32'b00010000001000000000000000000000;
          10'd512: delta_out = 32'b00010000000000000000000000000000;
          10'd513: delta_out = 32'b00001111111000000000000000000000;
        endcase
     end
endmodule
